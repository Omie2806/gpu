module imm_gen (
    input  logic [15:0] imm,      
    output logic [15:0] imm_out
);

    assign imm_out = imm;   

endmodule